library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_sprite_ram is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(8 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_sprite_ram is
	type rom is array(0 to  511) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"4F",X"B4",X"BC",X"00",X"4F",X"B4",X"B4",X"00",X"4F",X"6A",X"AC",X"00", -- modified
		X"4C",X"AA",X"81",X"00",X"00",X"00",X"B4",X"00",X"00",X"00",X"8C",X"00",X"00",X"00",X"80",X"00", -- modified		
--		X"00",X"00",X"00",X"00",X"4F",X"B4",X"BC",X"00",X"4F",X"B4",X"B4",X"00",X"4F",X"2A",X"AC",X"00", -- ori
--		X"4C",X"2A",X"81",X"00",X"00",X"00",X"B4",X"00",X"00",X"00",X"8C",X"00",X"00",X"00",X"80",X"00", -- ori
		X"00",X"00",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4A",X"07",X"C1",X"00", 
		X"47",X"06",X"D1",X"00",X"57",X"12",X"D1",X"00",X"47",X"16",X"E1",X"00",X"57",X"1A",X"E1",X"00", 
		X"45",X"00",X"C4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"36",X"29",X"23",X"00",X"36",X"29",X"30",X"00",X"36",X"2E",X"3D",X"00",X"4C",X"29",X"23",X"00",
		X"4C",X"29",X"30",X"00",X"4C",X"00",X"3D",X"00",X"62",X"29",X"23",X"00",X"62",X"2E",X"30",X"00",
		X"62",X"00",X"3D",X"00",X"78",X"2E",X"23",X"00",X"78",X"00",X"30",X"00",X"78",X"00",X"3D",X"00",
		X"8E",X"68",X"23",X"00",X"8E",X"00",X"30",X"00",X"8E",X"00",X"3D",X"00",X"A4",X"29",X"23",X"00",
		X"A4",X"29",X"30",X"00",X"A4",X"00",X"3D",X"00",X"BA",X"29",X"23",X"00",X"BA",X"2A",X"30",X"00",
		X"BA",X"2A",X"3D",X"00",X"D0",X"29",X"23",X"00",X"D0",X"2E",X"30",X"00",X"D0",X"29",X"3D",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"32",X"00",
		X"00",X"00",X"38",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"38",X"00",
		X"00",X"00",X"38",X"00",X"00",X"00",X"38",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"BE",X"B8",X"00",X"00",X"B9",X"B8",X"00",X"EC",X"2E",X"CA",X"00",X"EC",X"2A",X"B2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
