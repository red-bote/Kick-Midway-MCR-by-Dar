library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity kick_video_ram is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(9 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of kick_video_ram is
	type rom is array(0 to  1023) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"0E",X"14",X"12",X"0E",X"14",X"12",X"0E",X"14",X"12",X"0E",X"14",X"12",X"0E",X"14",X"12",X"0E",
		X"14",X"12",X"0E",X"14",X"12",X"0E",X"14",X"12",X"0E",X"14",X"12",X"0E",X"0B",X"14",X"14",X"12",
		X"0E",X"14",X"11",X"0E",X"14",X"11",X"0E",X"14",X"11",X"0E",X"14",X"11",X"0E",X"14",X"11",X"0E",
		X"14",X"11",X"0E",X"14",X"11",X"0E",X"14",X"11",X"0E",X"14",X"11",X"0E",X"0B",X"14",X"14",X"11",
		X"0D",X"15",X"10",X"0D",X"15",X"10",X"0D",X"15",X"10",X"0D",X"15",X"10",X"0D",X"15",X"10",X"0D",
		X"15",X"10",X"0D",X"15",X"10",X"0D",X"15",X"10",X"0D",X"15",X"10",X"0D",X"0A",X"15",X"15",X"10",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"5C",X"5F",X"5C",X"5F",
		X"5C",X"5F",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"D0",X"D0",X"D0",X"43",X"D0",X"D0",
		X"76",X"14",X"50",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"BB",X"5F",X"13",X"5F",
		X"13",X"5F",X"13",X"5F",X"13",X"13",X"13",X"13",X"BD",X"BC",X"D0",X"D0",X"D0",X"52",X"43",X"D0",
		X"14",X"14",X"4C",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"BF",X"5C",
		X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"5C",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"45",X"41",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"1C",X"C5",X"C4",X"91",
		X"91",X"91",X"91",X"91",X"5B",X"C3",X"C2",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"44",X"54",X"D0",
		X"14",X"14",X"31",X"30",X"14",X"14",X"14",X"14",X"14",X"23",X"1F",X"26",X"22",X"C6",X"C7",X"C8",
		X"C8",X"C8",X"C8",X"C8",X"C8",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"49",X"43",X"D0",
		X"14",X"14",X"76",X"14",X"14",X"14",X"14",X"14",X"14",X"1B",X"1B",X"22",X"22",X"22",X"E2",X"C6",
		X"C7",X"C8",X"C9",X"CA",X"CB",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"54",X"48",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"1F",X"22",X"26",X"22",X"22",X"22",
		X"14",X"14",X"14",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"53",X"D0",X"D0",
		X"14",X"14",X"48",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"1D",X"14",X"14",X"BA",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"42",X"D0",
		X"76",X"14",X"49",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"11",X"22",X"22",X"14",
		X"14",X"14",X"AA",X"B9",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"41",X"D0",
		X"14",X"14",X"14",X"32",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"1F",X"22",X"26",X"22",
		X"14",X"C8",X"CB",X"DE",X"B6",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"30",X"4C",X"D0",
		X"14",X"76",X"53",X"30",X"14",X"20",X"1E",X"26",X"22",X"22",X"26",X"22",X"22",X"22",X"22",X"14",
		X"B2",X"B3",X"A5",X"DF",X"DC",X"B4",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"4C",X"D0",
		X"14",X"14",X"43",X"30",X"14",X"14",X"20",X"1B",X"1B",X"1B",X"1E",X"22",X"26",X"22",X"22",X"E2",
		X"14",X"14",X"B0",X"DA",X"DF",X"B1",X"AD",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"4F",X"D0",
		X"14",X"14",X"4F",X"30",X"14",X"14",X"14",X"14",X"14",X"14",X"20",X"1B",X"1B",X"1B",X"1B",X"1E",
		X"14",X"AA",X"AB",X"DF",X"DC",X"DC",X"A9",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"4F",X"D0",
		X"14",X"14",X"52",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"22",X"E2",X"11",
		X"A7",X"A8",X"A8",X"DE",X"DC",X"DB",X"DA",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"4E",X"D0",
		X"14",X"14",X"45",X"14",X"14",X"14",X"14",X"14",X"14",X"1F",X"26",X"22",X"26",X"22",X"A6",X"9F",
		X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"9F",X"A2",X"A1",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"14",X"14",X"14",X"76",X"14",X"14",X"14",X"14",X"07",X"22",X"22",X"22",X"22",X"14",X"9E",X"99",
		X"9F",X"9F",X"5B",X"9F",X"9F",X"5C",X"9F",X"9F",X"A0",X"D0",X"D0",X"D0",X"D0",X"D0",X"4F",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"1C",X"E2",X"E2",X"9C",X"9A",X"9B",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"9D",X"D0",X"D0",X"D0",X"D0",X"4E",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"96",X"5B",X"91",X"91",X"91",X"91",
		X"91",X"5B",X"5B",X"5B",X"5B",X"91",X"91",X"5B",X"5B",X"CF",X"97",X"D0",X"D0",X"D0",X"D0",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"95",X"5B",X"91",X"91",X"5B",X"91",X"91",
		X"91",X"5B",X"91",X"91",X"91",X"91",X"5B",X"5B",X"5B",X"5B",X"98",X"D0",X"D0",X"D0",X"48",X"D0",
		X"14",X"76",X"14",X"14",X"14",X"14",X"14",X"14",X"90",X"91",X"91",X"91",X"92",X"93",X"93",X"93",
		X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"94",X"D0",X"D0",X"45",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"76",X"14",X"14",X"61",X"5C",X"5C",X"1A",X"13",X"13",X"5F",X"13",
		X"5F",X"13",X"5F",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"27",X"D0",X"D0",X"41",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"61",X"5C",X"5C",X"63",X"13",X"13",X"A4",X"13",
		X"A4",X"13",X"A4",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"D0",X"D0",X"44",X"D0",
		X"14",X"14",X"14",X"14",X"14",X"5D",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"5F",X"D0",X"D0",X"D0",X"D0",
		X"76",X"14",X"76",X"14",X"14",X"03",X"5C",X"06",X"03",X"5C",X"06",X"03",X"5C",X"06",X"03",X"5C",
		X"06",X"03",X"5C",X"06",X"03",X"5C",X"06",X"03",X"5C",X"06",X"03",X"5C",X"D0",X"D0",X"D0",X"D0",
		X"14",X"14",X"02",X"05",X"04",X"02",X"05",X"04",X"02",X"05",X"04",X"02",X"05",X"04",X"02",X"05",
		X"04",X"02",X"05",X"04",X"02",X"05",X"04",X"02",X"05",X"04",X"02",X"02",X"02",X"02",X"02",X"02",
		X"14",X"14",X"09",X"07",X"07",X"09",X"07",X"07",X"09",X"07",X"07",X"09",X"07",X"07",X"09",X"07",
		X"07",X"09",X"07",X"07",X"09",X"07",X"07",X"09",X"07",X"07",X"09",X"07",X"07",X"09",X"07",X"07",
		X"76",X"14",X"08",X"07",X"07",X"08",X"07",X"07",X"08",X"07",X"07",X"08",X"07",X"07",X"08",X"07",
		X"07",X"08",X"07",X"07",X"08",X"07",X"07",X"08",X"07",X"07",X"08",X"07",X"07",X"08",X"07",X"07",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",
		X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14",X"14");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
